use ieee;
